module top(
    //ports
    input bit clock,
    input bit reset,
    //outport
);

//wire declarations
//regs declarations

//logic blocks

endmodule;
